/escnfs/courses/fa22-cse-40462.01/dropbox/dgarci23/mips8/muddlib.lef